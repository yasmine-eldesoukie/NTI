/*module edge_detector (
    input wire clk, rst,
    input wire in_signal,
    output reg edge
);

always @(posedge clk or negedge rst) begin
    if (!rst) begin
        
    end
end
endmodule
*/